module Lshift #(parameter WIDTH=32)(
  input [WIDTH-1:0] A,
  input [WIDTH-1:0] B,
  output [WIDTH-1:0] S
);
 wire [31:0] S0,S1,S2,S3;
    mux2 st0(S0, A, {A[30:0],1'b0},B[0]);
    mux2 st1(S1, S0, {S0[29:0],2'b0},B[1]);
    mux2 st2(S2, S1, {S1[27:0],4'b0},B[2]);
    mux2 st3(S3, S2, {S2[23:0],8'b0},B[3]);
    mux2 st4(S, S3, {S3[15:0],16'b0},B[4]);
endmodule



// module Lshift #(parameter WIDTH=32)(
//   input [WIDTH-1:0] data_in,       
//     input [5:0] shift_amount,   
//     input load,                 
//   output reg [WIDTH-1:0] data_out  
// );

//   reg [WIDTH-1:0] shifted_data;  
// integer i;
// always @* begin
//     if (load) begin
//         shifted_data = data_in;
//         for (i = 0; i < shift_amount; i = i + 1) begin
//             shifted_data = {shifted_data[30:0], 1'b0}; 
//         end
//     end
// end

// always @* begin
//     data_out = shifted_data;
// end

// endmodule
